// Code your design here
// F = (A'+B'+C).(A'+B'+C').(A+B+C).(A+B+C'), dataflow

module sop(a,b,c,y);

input a,b,c;
output y;
assign y = (~a|~b|c)&(~a|~b|~c)&(a|b|c)&(a|b|~c);

endmodule
